module Equal (in_equal, out_equal);
  input [31:0] in_equal;
  output out_equal;
  
  or or0_0(out_equal, in_equal[0], in_equal[1], in_equal[2], in_equal[3], in_equal[4], in_equal[5], in_equal[6], in_equal[7], in_equal[8], in_equal[9], in_equal[10], in_equal[11], in_equal[12], in_equal[13], in_equal[14], in_equal[15], in_equal[16], in_equal[17], in_equal[18], in_equal[19], in_equal[20], in_equal[21], in_equal[22], in_equal[23], in_equal[24], in_equal[25], in_equal[26], in_equal[27], in_equal[28], in_equal[29], in_equal[30], in_equal[31]);
endmodule
