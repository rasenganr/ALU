module myNOT (in_not, out_not);
  input [31:0] in_not;
  output [31 :0] out_not;
  
  not not0(out_not[0], in_not[0]);
  not not1(out_not[1], in_not[1]);
  not not2(out_not[2], in_not[2]);
  not not3(out_not[3], in_not[3]);
  not not4(out_not[4], in_not[4]);
  not not5(out_not[5], in_not[5]);
  not not6(out_not[6], in_not[6]);
  not not7(out_not[7], in_not[7]);
  not not8(out_not[8], in_not[8]);
  not not9(out_not[9], in_not[9]);
  not not10(out_not[10], in_not[10]);
  not not11(out_not[11], in_not[11]);
  not not12(out_not[12], in_not[12]);
  not not13(out_not[13], in_not[13]);
  not not14(out_not[14], in_not[14]);
  not not15(out_not[15], in_not[15]);
  not not16(out_not[16], in_not[16]);
  not not17(out_not[17], in_not[17]);
  not not18(out_not[18], in_not[18]);
  not not19(out_not[19], in_not[19]);
  not not20(out_not[20], in_not[20]);
  not not21(out_not[21], in_not[21]);
  not not22(out_not[22], in_not[22]);
  not not23(out_not[23], in_not[23]);
  not not24(out_not[24], in_not[24]);
  not not25(out_not[25], in_not[25]);
  not not26(out_not[26], in_not[26]);
  not not27(out_not[27], in_not[27]);
  not not28(out_not[28], in_not[28]);
  not not29(out_not[29], in_not[29]);
  not not30(out_not[30], in_not[30]);
  not not31(out_not[31], in_not[31]);
endmodule
